library verilog;
use verilog.vl_types.all;
entity mips_core is
    port(
        clock           : in     vl_logic
    );
end mips_core;
